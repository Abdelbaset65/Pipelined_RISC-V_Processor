

module singleMem (input         clk, s_clk,
                                MemRead,
                                MemWrite,
                  input  [2:0]  func,
                  input  [5:0]  addr,
                  input  [31:0] data_in,
                  output reg [31:0] data_out);


    reg [7:0] mem [0:511];
    always@(posedge s_clk)begin
    data_out = mem[addr];
    end
    always@(negedge clk)begin
    data_out =  MemRead ? {mem[addr+255], mem[addr+255+1], mem[addr+255+2], mem[addr+255+3]}: 0;
    end
    initial 
    begin
        mem[255]=8'd25;
        mem[256]=8'd25;
    end 

    always @(posedge clk)begin
    if(MemWrite)
    case(func)
    3'b000:mem[addr+255] <= data_in[7:0];
    3'b001:{mem[addr+255], mem[addr+255+1]} <= data_in[15:0];
    3'b010:{mem[addr+255], mem[addr+255+1], mem[addr+255+2], mem[addr+255+3]} <= data_in;
    endcase 
    end

    initial 
    begin
      {mem[3],  mem[2],  mem[1],  mem[0]}  = 32'b00000000000000000011000100010111;
      {mem[7],  mem[6],  mem[5],  mem[4]}  = 32'b00000000000000001100000010110111;
      {mem[11], mem[10], mem[9],  mem[8]}  = 32'b00000010000000000000000111101111;
      {mem[15], mem[14], mem[13], mem[12]} = 32'b00000000010000010000000111100111;
      {mem[19], mem[18], mem[17], mem[16]} = 32'b00000000000100010000010001100011;
      {mem[23], mem[22], mem[21], mem[20]} = 32'b00000000000100010001001001100011;
      {mem[27], mem[26], mem[25], mem[24]} = 32'b00000000000100010100100001100011;
      {mem[31], mem[30], mem[29], mem[28]} = 32'b00000000000100010101011001100011;
      {mem[35], mem[34], mem[33], mem[32]} = 32'b00000000100000010000000100000011;
      {mem[39], mem[38], mem[37], mem[36]} = 32'b00000001000000010010000100000011;
      {mem[43], mem[42], mem[41], mem[40]} = 32'b00000000000100010000001000100011;
      {mem[47], mem[46], mem[45], mem[44]} = 32'b00000000000100010010100000100011;
      {mem[51], mem[50], mem[49], mem[48]} = 32'b00000001000000001100000100000011;
      {mem[55], mem[54], mem[53], mem[52]} = 32'b00000001010000010000000110010011;
      {mem[59], mem[58], mem[57], mem[56]} = 32'b00000000001000011010000110010011;
      {mem[63], mem[62], mem[61], mem[60]} = 32'b11111111111000011011000110010011;
      {mem[67], mem[66], mem[65], mem[64]} = 32'b00000001111000011100000110010011;
      {mem[71], mem[70], mem[69], mem[68]} = 32'b00000000000100011111001000110011;
      {mem[75], mem[74], mem[73], mem[72]} = 32'b00000000001100100000001010110011;
      {mem[79], mem[78], mem[77], mem[76]} = 32'b00000000000000000000000001110011;
      {mem[83], mem[82], mem[81], mem[80]} = 32'b00000000000100000000000001110011;
      {mem[87], mem[86], mem[85], mem[84]} = 32'b01000000001000101101001100110011;
      {mem[91], mem[90], mem[89], mem[88]} = 32'b00000000000100110010001110110011;
      {mem[95], mem[94], mem[93], mem[92]} = 32'b11111010001000011111111011100011;
    end

endmodule