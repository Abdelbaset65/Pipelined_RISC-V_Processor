`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/06/2020 09:12:40 AM
// Design Name: 
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////




module InstMem (input [5:0] addr, output [31:0] data_out);
 reg [31:0] mem [0:63];
 assign data_out = mem[addr];

initial begin
//mem[0]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//mem[1]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
//mem[2]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
//mem[3]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
//mem[4]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
//mem[5]=32'b0_000000_00011_00100_000_0100_0_1100011 ; //beq x4, x3, L
//mem[6]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
//mem[7]=32'b0000000_00010_00011_000_00101_0110011 ; //L: add x5,x3,x2
//mem[8]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
//mem[9]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
//mem[10]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
//mem[11]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
//mem[12]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
//mem[13]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1

mem[0]=32'b00000000000001100100000010110111
mem[1]=32'b00000000000000010100000100010111
mem[2]=32'b00000000100000010000000111100111
mem[3]=32'b00000000010000000000010011101111
mem[4]=32'b00000000001100010000111001100011
mem[5]=32'b00000000001100010001110001100011
mem[6]=32'b00000000001100010100101001100011
mem[7]=32'b00000000001100010101100001100011
mem[8]=32'b00000000001100010110011001100011
mem[9]=32'b00000000001100010111010001100011
mem[10]=32'b00000001010000011000000100000011
mem[11]=32'b00000000001000011001000100000011
mem[12]=32'b00000000010000011010000100000011
mem[13]=32'b00000000100000011100000100000011
mem[14]=32'b00000000110000011101000100000011
mem[15]=32'b00000000001000011000010100100011
mem[16]=32'b00000000001000011001011000100011
mem[17]=32'b00000000001000011010011000100011
mem[18]=32'b00000000101000011000000100010011
mem[19]=32'b11111111011000011010000100010011
mem[20]=32'b11111111011000011011000100010011
mem[21]=32'b00111110100000011100001000010011
mem[22]=32'b00000001100100011111001000010011
mem[23]=32'b00000001100100011001001010010011
mem[24]=32'b00000000011100011101001100010011
mem[25]=32'b01000000011000100101000110010011
mem[26]=32'b00000000001000011000001000110011
mem[27]=32'b01000000001100100000000100110011
mem[28]=32'b00000000010100101001001100110011
mem[29]=32'b00000000001000011010001010110011
mem[30]=32'b00000000001000011011001010110011
mem[31]=32'b00000000001000011100001000110011
mem[32]=32'b00000000000100011101001110110011
mem[33]=32'b01000000000000001101000100110011
mem[34]=32'b00000000010100011110000010110011
mem[35]=32'b00000000011000111111000100110011
mem[36]=32'b00000000000000000000000001110011
mem[37]=32'b00000000000100000000000001110011





// mem[0]= 32'b00000000000000000010000010000011; //lw x1, 0(x0)
// mem[1]= 32'b00000000010000000010000100000011; //lw x2, 4(x0)
// mem[2]= 32'b00000000001000001000000110110011; //add x3, x1, x2
// mem[3]= 32'b01000000001000001000001000110011; //sub x4, x1, x2
// mem[4]= 32'b00000000001000001111001010110011; //and x5, x1, x2
// mem[5]= 32'b00000000001000001110001100110011; //or x6, x1, x2
// mem[6]= 32'b00000000000000100000010001100011; //beq x4, x0, L1
// mem[7]= 32'b00000000010000000010010000100011; //sw x4, 8(x0)
// mem[8]= 32'b00000000001100000010010000100011; //L1: sw x3, 8(x0)                                               
end

endmodule